// `timescale 1ns / 1ps

// module Mult(
//             input 

//     );
// endmodule
